netcdf PLDP_1km_nc4_template {
dimensions:
	lon = 101 ;
	lat = 101 ;
	time = UNLIMITED ; // (0 currently)
variables:
	double time(time) ;
		time:longname = "Time" ;
		time:units = "days since 2001-01-01 00:00:00" ;
	float lon(lon) ;
		lon:longname = "Longitude" ;
		lon:shortname = "lon" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = -999.f ;
	float lat(lat) ;
		lat:longname = "Latitude" ;
		lat:shortname = "lat" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = -999.f ;
	float u(time, lat, lon) ;
		u:longname = "Eastward Velocity" ;
		u:standard_name = "eastward_surface_velocity" ;
		u:shortname = "u" ;
		u:units = "cm/s" ;
		u:_FillValue = -999.f ;
	float v(time, lat, lon) ;
		v:longname = "Northward Velocity" ;
		v:standard_name = "northward_surface_velocity" ;
		v:shortname = "v" ;
		v:units = "cm/s" ;
		v:_FillValue = -999.f ;
	float u_err(time, lat, lon) ;
		u_err:_FillValue = -999.f ;
	float v_err(time, lat, lon) ;
		v_err:_FillValue = -999.f ;
	int num_radials(time, lat, lon) ;
		num_radials:_FillValue = -999 ;
	int site_code(time, lat, lon) ;
		site_code:_FillValue = -999 ;

// global attributes:
		:history = "Converted into netCDF by process_codar_totals_into_netcdf" ;
		:source = "/Users/codar/Desktop/Data/PLDP/oi/ascii/*" ;
		:header = "\n",
			"%TimeStamp: 2009 01 01 00 00\n",
			"%TimeZone: GMT+0.000\n",
			"%Domain: BPU\n",
			"%Type: OI\n",
			"%DataCreationInfo: Rutgers/BPU Domain\n",
			"%DataCreationTimeStamp: 01-Apr-2009 23:12:51\n",
			"%DataCreationTimeZone: GMT\n",
			"%ProcessingProgram: TUVstruct2ascii_OI 06-Apr-2009 17:54:14\n",
			"%TUV_structVersion: SVN $Rev: 396 $ $Date: 2007-04-02 16:56:29 +0000 (Mon, 02 Apr 2007) $\n",
			"%MinNumSites:    2\n",
			"%MinNumRads:   3\n",
			"%mdlvar: 420.00\n",
			"%errvar:  66.00\n",
			"%sx:  5.00\n",
			"%sy:  8.00\n",
			"%tempthresh: 0.020833\n";
			
			data:
			
			lon = -65.501906, -65.480991, -65.460077, -65.439162, -65.418247, -65.397332, -65.376418, -65.355503, -65.334588, -65.313673, -65.292759, -65.271844, -65.250929, -65.230014, -65.209100, -65.188185, -65.167270, -65.146355, -65.125441, -65.104526, -65.083611, -65.062696, -65.041782, -65.020867, -64.999952, -64.979038, -64.958123, -64.937208, -64.916293, -64.895379, -64.874464, -64.853549, -64.832634, -64.811720, -64.790805, -64.769890, -64.748975, -64.728061, -64.707146, -64.686231, -64.665316, -64.644402, -64.623487, -64.602572, -64.581657, -64.560743, -64.539828, -64.518913, -64.497998, -64.477084, -64.456169, -64.435254, -64.414340, -64.393425, -64.372510, -64.351595, -64.330681, -64.309766, -64.288851, -64.267936, -64.247022, -64.226107, -64.205192, -64.184277, -64.163363, -64.142448, -64.121533, -64.100618, -64.079704, -64.058789, -64.037874, -64.016959, -63.996045, -63.975130, -63.954215, -63.933301, -63.912386, -63.891471, -63.870556, -63.849642, -63.828727, -63.807812, -63.786897, -63.765983, -63.745068, -63.724153, -63.703238, -63.682324, -63.661409, -63.640494, -63.619579, -63.598665, -63.577750, -63.556835, -63.535920, -63.515006, -63.494091, -63.473176, -63.452261, -63.431347, -63.410432;
			
			lat = -65.432216, -65.423223, -65.414230, -65.405236, -65.396243, -65.387250, -65.378257, -65.369264, -65.360270, -65.351277, -65.342284, -65.333291, -65.324297, -65.315304, -65.306311, -65.297318, -65.288325, -65.279331, -65.270338, -65.261345, -65.252352, -65.243359, -65.234365, -65.225372, -65.216379, -65.207386, -65.198393, -65.189399, -65.180406, -65.171413, -65.162420, -65.153426, -65.144433, -65.135440, -65.126447, -65.117454, -65.108460, -65.099467, -65.090474, -65.081481, -65.072488, -65.063494, -65.054501, -65.045508, -65.036515, -65.027522, -65.018528, -65.009535, -65.000542, -64.991549, -64.982555, -64.973562, -64.964569, -64.955576, -64.946583, -64.937589, -64.928596, -64.919603, -64.910610, -64.901617, -64.892623, -64.883630, -64.874637, -64.865644, -64.856651, -64.847657, -64.838664, -64.829671, -64.820678, -64.811685, -64.802691, -64.793698, -64.784705, -64.775712, -64.766718, -64.757725, -64.748732, -64.739739, -64.730746, -64.721752, -64.712759, -64.703766, -64.694773, -64.685780, -64.676786, -64.667793, -64.658800, -64.649807, -64.640814, -64.631820, -64.622827, -64.613834, -64.604841, -64.595847, -64.586854, -64.577861, -64.568868, -64.559875, -64.550881, -64.541888, -64.532895;
			
}

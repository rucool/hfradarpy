netcdf NY_1km_nc4_template {
dimensions:
	lon = 79 ;
	lat = 45 ;
	time = UNLIMITED ; // (0 currently)
variables:
	double time(time) ;
		time:longname = "Time" ;
		time:units = "days since 2001-01-01 00:00:00" ;
	float lon(lon) ;
		lon:longname = "Longitude" ;
		lon:shortname = "lon" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = -999.f ;
	float lat(lat) ;
		lat:longname = "Latitude" ;
		lat:shortname = "lat" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = -999.f ;
	float u(time, lat, lon) ;
		u:longname = "Eastward Velocity" ;
		u:standard_name = "eastward_surface_velocity" ;
		u:shortname = "u" ;
		u:units = "cm/s" ;
		u:_FillValue = -999.f ;
	float v(time, lat, lon) ;
		v:longname = "Northward Velocity" ;
		v:standard_name = "northward_surface_velocity" ;
		v:shortname = "v" ;
		v:units = "cm/s" ;
		v:_FillValue = -999.f ;
	float u_err(time, lat, lon) ;
		u_err:_FillValue = -999.f ;
	float v_err(time, lat, lon) ;
		v_err:_FillValue = -999.f ;
	int num_radials(time, lat, lon) ;
		num_radials:_FillValue = -999 ;
	int site_code(time, lat, lon) ;
		site_code:_FillValue = -999 ;

// global attributes:
		:history = "Converted into netCDF by process_codar_totals_into_netcdf" ;
		:source = "/Users/codar/Desktop/Data/mara/oi/ascii/*" ;
		:header = "\n",
			"%TimeStamp: 2009 01 01 00 00\n",
			"%TimeZone: GMT+0.000\n",
			"%Domain: NYH\n",
			"%Type: OI\n",
			"%DataCreationInfo: Rutgers/NYH Domain\n",
			"%DataCreationTimeStamp: 01-Apr-2009 23:12:51\n",
			"%DataCreationTimeZone: GMT\n",
			"%ProcessingProgram: TUVstruct2ascii_OI 06-Apr-2009 17:54:14\n",
			"%TUV_structVersion: SVN $Rev: 396 $ $Date: 2007-04-02 16:56:29 +0000 (Mon, 02 Apr 2007) $\n",
			"%MinNumSites:    2\n",
			"%MinNumRads:   3\n",
			"%mdlvar: 420.00\n",
			"%errvar:  66.00\n",
			"%sx:  5.00\n",
			"%sy:  8.00\n",
			"%tempthresh: 0.020833\n";
			
			data: 
			
			lon = -74.256922, -74.247243, -74.237564, -74.227884, -74.218205, -74.208526, -74.198847, -74.189168, -74.179488, -74.169809, -74.160130, -74.150451, -74.140772, -74.131093, -74.121413, -74.111734, -74.102055, -74.092376, -74.082697, -74.073017, -74.063338, -74.053659, -74.043980, -74.034301, -74.024621, -74.014942, -74.005263, -73.995584, -73.985905, -73.976225, -73.966546, -73.956867, -73.947188, -73.937509, -73.927829, -73.918150, -73.908471, -73.898792, -73.889113, -73.879434, -73.869754, -73.860075, -73.850396, -73.840717, -73.831038, -73.821358, -73.811679, -73.802000, -73.792321, -73.782642, -73.772962, -73.763283, -73.753604, -73.743925, -73.734246, -73.724566, -73.714887, -73.705208, -73.695529, -73.685850, -73.676170, -73.666491, -73.656812, -73.647133, -73.637454, -73.627775, -73.618095, -73.608416, -73.598737, -73.589058, -73.579379, -73.569699, -73.560020, -73.550341, -73.540662, -73.530983, -73.521303, -73.511624, -73.501945;
			
			lat = 40.201420, 40.210410, 40.219400, 40.228390, 40.237380, 40.246370, 40.255360, 40.264350, 40.273340, 40.282330, 40.291320, 40.300310, 40.309300, 40.318290, 40.327280, 40.336270, 40.345260, 40.354250, 40.363240, 40.372230, 40.381220, 40.390210, 40.399200, 40.408190, 40.417180, 40.426170, 40.435160, 40.444150, 40.453140, 40.462130, 40.471120, 40.480110, 40.489100, 40.498090, 40.507080, 40.516070, 40.525060, 40.534050, 40.543040, 40.552030, 40.561020, 40.570010, 40.579000, 40.587990, 40.596980;
			
}
